//1.definicion del modulo y sus I/O
//Dentro del parentesis se define los I/O

module _and( input a,input b, output c );
//2.Define cables o componentes internos
//NA
//3.Asignaciones,Instancias y conexiones

assign c = a & b;

endmodule
